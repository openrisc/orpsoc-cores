`include "timescale.v"

module orpsoc_tb;

   vlog_tb_utils vlog_tb_utils0();

   ////////////////////////////////////////////////////////////////////////
   //
   // ELF program loading
   // 
   ////////////////////////////////////////////////////////////////////////
   integer mem_words;
   integer i;
   reg [31:0] mem_word;
   reg [1023:0] elf_file;

   initial begin
      if($value$plusargs("elf_load=%s", elf_file)) begin
	 $elf_load_file(elf_file);
	 
	 mem_words = $elf_get_size/4;
	 $display("Loading %d words", mem_words);
	 for(i=0; i < mem_words; i = i+1)
	   orpsoc_tb.dut.wb_bfm_memory0.mem[i] = $elf_read_32(i*4);
      end else
	$display("No ELF file specified");
      
   end

   ////////////////////////////////////////////////////////////////////////
   //
   // Clock and reset generation
   // 
   ////////////////////////////////////////////////////////////////////////
   reg wb_clk = 1;
   reg wb_rst = 1;

   always #5 wb_clk <= ~wb_clk;
   initial #100 wb_rst <= 0;

   ////////////////////////////////////////////////////////////////////////
   //
   // OR1200 monitor
   // 
   ////////////////////////////////////////////////////////////////////////
   or1200_monitor i_monitor();
   
   ////////////////////////////////////////////////////////////////////////
   //
   // DUT
   // 
   ////////////////////////////////////////////////////////////////////////
   orpsoc_top
     #(.UART_SIM (1))
   dut
     (.wb_clk_i (wb_clk),
      .wb_rst_i (wb_rst));

endmodule
