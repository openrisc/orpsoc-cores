@00000000
00000013
20000093
00008067
	 
