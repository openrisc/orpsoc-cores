@00000000
18000000
18200000
A82104E2
BC010000
0FFFFFFF
9C21FFFF
18200000
A8210000
1880B000
A8400051
D8041000
D8040004
A8C00001
D8043004
04000018
A8600003
04000016
A8600000
04000014
A8600000
04000012
A8600000
18C00000
18E0FFFF
0400000E
E1013000
D8081800
9CC60001
BC060004
10000007
E4063800
0FFFFFF9
15000000
A8210100
44000800
D8040004
03FFFFF4
84E10000
D8041802
A8600001
A4630001
BC030001
13FFFFFE
8C640001
44004800
8C640002
	 
