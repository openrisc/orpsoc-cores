@00000000
18000000 A8200000 A8C00100 44003000
15000000 00000000 00000000 00000000
