//
// orpsoc-defines
//
`define MOR1KX
`ifndef MOR1KX
`define OR1200
`endif
`define UART0
`define SPI0
`define VGA0
`define ETH0
`define AC97
`define PS2_0
`define PS2_1
`define PS2_2
`define JTAG_DEBUG
`define RAM_WB
`define BOOTROM
// end of included module defines - keep this comment line here
